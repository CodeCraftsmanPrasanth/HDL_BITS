module top_module (
    input clk,
    input a,
    output q );
    always @(posedge clk) begin
        if(~a) q=1;
        else q=0;
    end
endmodule
